`include "uvm_macros.svh"
import uvm_pkg::*;

`include "seq_item.sv"
`include "sequencer.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "coverage.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
`include "wr_test.sv"
`include "rd_test.sv"
`include "wr_rd_test.sv"
`include "wr_rd_low_test.sv"
`include "wr_after_rd_test.sv"
`include "wr_rd_same_addr_test.sv"
`include "rd_only_particular_addr_test.sv"
`include "wr_rd_idle_test.sv"
`include "dut.sv"
`include "interface.sv"
`include "testbench.sv"



